`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NetWalk
// Engineer: Mahesh Dananjaya
// 
// Create Date: 01/07/2016 03:15:47 PM
// Design Name: 
// Module Name: netwalk_classification_engine
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module netwalk_classification_engine
#(parameter ADDR_WIDTH=32,PKT_BUFF_ADDR_WIDTH=9,OF_FLOW_TAG_WIDTH=5,DPL_PKT_BYTE_WIDTH=64,DPL_PKT_BIT_WIDTH=512,DPL_MATCH_FIELD_WIDTH=356, DPL_PKT_ADDR_WIDTH=6, DPL_PKT_DATA_WIDTH=8)
(
clk,
reset,

glbl_program_en,

pkt_header_ready,
pkt_header_accept,
//pkt_header_ready_accept,
//pkt_header_finish,
//pkt_header_finish_accept,
pkt_header_in,
pkt_header_data_buff,
sdn_match_field_ready,

//pkt_header_addr,
//pkt_header_data,
//pkt_header_read_enable,
/*
sdn_match_field_data,
sdn_match_field_ready,
sdn_match_field_accept,

sdn_ingress_port,
sdn_meta_data,
sdn_src_mac_addr,
sdn_dst_mac_addr,
sdn_ether_type,
sdn_vlan_id,
sdn_vlan_priority,
sdn_mpls_label,
sdn_mpls_fec_class,
sdn_src_ipv4_addr,
sdn_dst_ipv4_addr,
sdn_ipv4_protocol,
sdn_ipv4_tos,
sdn_tcp_src_port,
sdn_tcp_dst_port,
*/

OF_INGRESS_PORT,
OF_META_DATA,
OF_DST_MAC_ADDR,
OF_SRC_MAC_ADDR,
OF_ETHER_TYPE,
OF_VLAN_ID,
OF_VLAN_PRIORITY,
OF_MPLS_LABEL,
OF_MPLS_FEC_CLASS,
OF_SRC_IPV4_ADDR,
OF_DST_IPV4_ADDR,
OF_IP_PROTOCOL,
OF_IPV4_TOS,
OF_TCP_SRC_PORT,
OF_TCP_DST_PORT,

OF_MATCH_FIELD_DATA,
OF_FLOW_FOUND,

of_flow_tag,
openflow_packet_found,
packet_to_switch_found,

OF_INGRESS_PORT_ADDR,
OF_META_DATA_ADDR,
OF_DST_MAC_ADDR_ADDR,
OF_SRC_MAC_ADDR_ADDR,
OF_ETHER_TYPE_ADDR,
OF_VLAN_ID_ADDR,
OF_VLAN_PRIORITY_ADDR,
OF_MPLS_LABEL_ADDR,
OF_MPLS_FEC_CLASS_ADDR,
OF_SRC_IPV4_ADDR_ADDR,
OF_DST_IPV4_ADDR_ADDR,
OF_IP_PROTOCOL_ADDR,
OF_IPV4_TOS_ADDR,
OF_TCP_SRC_PORT_ADDR,
OF_TCP_DST_PORT_ADDR,

pkt_header_out,

pkt_addr_in,
pkt_addr_out

);

input [(ADDR_WIDTH*15)-1:0] pkt_addr_in;
output [(ADDR_WIDTH*15)-1:0] pkt_addr_out;

parameter INGRESS_PORT_WIDTH		=32;
parameter METADATA_WIDTH			=64;

parameter IP_ENCAP_WIDTH			=160;
parameter ETHER_ENCAP_WIDTH		=112;
parameter UDP_ENCAP_WIDTH			=64;
parameter TCP_ENCAP_WIDTH			=160;
parameter VLAN_ENCAP_WIDTH			=32;
parameter MPLS_ENCAP_WIDTH			=32;

//FIELD WIDTHS OF NETWORK STACK
parameter MAC_ADDR_WIDTH				=48;
parameter SRC_MAC_ADDR_WIDTH			=48;
parameter DST_MAC_ADDR_WIDTH			=48;
parameter ETHER_TYPE_WIDTH				=16;

parameter VLAN_TPID_WIDTH			=16;
parameter VLAN_PRIORITY_WIDTH		=3;
parameter VLAN_CFI_WIDTH			=1;
parameter VLAN_ID_WIDTH				=12;

parameter MPLS_LABEL_WIDTH			=20;
parameter MPLS_COS_WIDTH			=3;
parameter MPLS_S_WIDTH				=1;
parameter MPLS_TTL_WIDTH			=8;

parameter MPLS_FEC_WIDTH			=3;
parameter MPLS_FEC_CLASS_WIDTH			=3;

parameter IP_VERSION_WIDTH			=4;
parameter IP_IHL_WIDTH				=4;
parameter IP_DSCP_WIDTH				=6;
parameter IP_ECN_WIDTH				=2;
parameter IP_LENGTH_WIDTH			=16;
parameter IP_ID_WIDTH				=16;
parameter IP_FLAG_WIDTH				=3;
parameter IP_FRAGOFF_WIDTH			=13;
parameter IP_TTL_WIDTH				=8;
parameter IP_PROTOCOL_WIDTH		=8;
parameter IP_CHECKSUM_WIDTH		=16;
parameter IP_ADDR_WIDTH				=32;
parameter IP_SRC_ADDR_WIDTH				=32;
parameter IP_DST_ADDR_WIDTH				=32;

//parameter IP_TOS_WIDTH=IP_DSCP_WIDTH+IP_ECN_WIDTH;
parameter IP_TOS_WIDTH=IP_DSCP_WIDTH;

parameter TCP_PORT_WIDTH			=16;
parameter TCP_SRC_PORT_WIDTH		=16;
parameter TCP_DST_PORT_WIDTH		=16;
parameter TCP_SEQN_WIDTH			=32;
parameter TCP_ACKN_WIDTH			=32;
parameter TCP_DTOFF_WIDTH			=4;
parameter TCP_RESV_WIDTH			=3;
parameter TCP_NS_WIDTH				=1;
parameter TCP_CWR_WIDTH				=1;
parameter TCP_ECE_WIDTH				=1;
parameter TCP_UGR_WIDTH				=1;
parameter TCP_ACK_WIDTH				=1;
parameter TCP_PSH_WIDTH				=1;
parameter TCP_RST_WIDTH				=1;
parameter TCP_SYN_WIDTH				=1;
parameter TCP_FIN_WIDTH				=1;
parameter TCP_WINSIZE_WIDTH		=16;
parameter TCP_CHECKSUM_WIDTH		=16;
parameter TCP_URGPNT_WIDTH			=16;

parameter UDP_PORT_WIDTH			=16;
parameter UDP_SRC_PORT_WIDTH		=16;
parameter UDP_DST_PORT_WIDTH		=16;
parameter UDP_LENGTH_WIDTH			=16;
parameter UDP_CHECKSUM_WIDTH		=16;

//FIELD OFFSET
parameter INGRESS_PORT_OFFSET   =0;
parameter METADATA_OFFSET		  =32;

parameter MAC_DST_OFFSET			=0;
parameter MAC_SRC_OFFSET			=MAC_ADDR_WIDTH;
parameter ETHER_TYPE_OFFSET		=MAC_ADDR_WIDTH+MAC_ADDR_WIDTH;

parameter VLAN_TPID_OFFSET			=0;
parameter VLAN_PRIORITY_OFFSET	=16;
parameter VLAN_CFI_OFFSET			=19;
parameter VLAN_ID_OFFSET			=20;

parameter MPLS_LABEL_OFFSET		=0;
parameter MPLS_COS_OFFSET			=20;
parameter MPLS_S_OFFSET				=23;
parameter MPLS_TTL_OFFSET			=24;
parameter MPLS_FEC_OFFSET			=20;
parameter MPLS_FEC_CLASS_OFFSET	=3;

parameter IP_VERSION_OFFSET		=0;
parameter IP_IHL_OFFSET				=4;
parameter IP_DSCP_OFFSET			=8;
parameter IP_ECN_OFFSET				=14;
parameter IP_LENGTH_OFFSET			=16;
parameter IP_ID_OFFSET				=32;
parameter IP_FLAG_OFFSET			=48;
parameter IP_FRAGOFF_OFFSET			=51;
parameter IP_TTL_OFFSET				=64;
parameter IP_PROTOCOL_OFFSET		=72;
parameter IP_CHECKSUM_OFFSET		=80;
parameter IP_SRC_ADDR_OFFSET		=96;
parameter IP_DST_ADDR_OFFSET		=128;
parameter IP_TOS_OFFSET				=8;

parameter TCP_SRC_PORT_OFFSET			=0;
parameter TCP_DST_PORT_OFFSET			=16;
parameter TCP_SEQN_OFFSET			=32;
parameter TCP_ACKN_OFFSET			=64;
parameter TCP_DTOFF_OFFSET			=96;
parameter TCP_RESV_OFFSET			=100;
parameter TCP_NS_OFFSET				=103;
parameter TCP_CWR_OFFSET				=104;
parameter TCP_ECE_OFFSET				=105;
parameter TCP_UGR_OFFSET				=106;
parameter TCP_ACK_OFFSET				=107;
parameter TCP_PSH_OFFSET				=108;
parameter TCP_RST_OFFSET				=109;
parameter TCP_SYN_OFFSET				=110;
parameter TCP_FIN_OFFSET				=111;
parameter TCP_WINSIZE_OFFSET		=112;
parameter TCP_CHECKSUM_OFFSET		=128;
parameter TCP_URGPNT_OFFSET			=142;

parameter UDP_SRC_PORT_OFFSET			=0;
parameter UDP_DST_PORT_OFFSET			=16;
parameter UDP_LENGTH_OFFSET			=32;
parameter UDP_CHECKSUM_OFFSET		   =48;

//TREE CLASSIFICATION PATHS
parameter ROOT_ADDR									=0;
parameter BASE_ADDR									=96;//32;   //BASE ADDRESS
parameter ETHER_HEAD									=BASE_ADDR;
parameter ETHER_ARP_HEAD							=BASE_ADDR+ETHER_ENCAP_WIDTH;
//parameter ETHER_VLAN_ETHER_HEAD		=BASE_ADDR;
parameter ETHER_VLAN_FLOW_VLAN_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH;

parameter ETHER_VLAN_ARP_FLOW_VLAN_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_ARP_FLOW_ARP_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;

parameter ETHER_MPLS_FLOW_MPLS_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH;

parameter ETHER_IP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH;

parameter ETHER_VLAN_MPLS_FLOW_VLAN_HEAD		=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_FLOW_MPLS_HEADER	=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;

parameter ETHER_VLAN_IP_FLOW_VLAN_HEAD 		=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_FLOW_IP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;

parameter ETHER_MPLS_IP_FLOW_MPLS_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_FLOW_IP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;

parameter ETHER_IP_TCP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_IP_TCP_FLOW_TCP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_IP_UDP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_IP_UDP_FLOW_UDP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+IP_ENCAP_WIDTH;

//OPTIONAL
parameter ETHER_IP_ICMP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_IP_ICMP_FLOW_ICMP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+IP_ENCAP_WIDTH;
//OPTIONAL

parameter ETHER_VLAN_MPLS_IP_FLOW_VLAN_HEAD		   	=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_FLOW_MPLS_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;

parameter ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD 		=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_TCP_FLOW_IP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD 		=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_UDP_FLOW_IP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD 		=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_IP_ICMP_FLOW_ICMP_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_TCP_FLOW_IP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_UDP_FLOW_IP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD			=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_MPLS_IP_ICMP_FLOW_ICMP_HEAD			   =BASE_ADDR+ETHER_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD		   	=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD		   	=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

parameter ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD		   	=BASE_ADDR+ETHER_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD				=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH;
parameter ETHER_VLAN_MPLS_IP_ICMP_FLOW_ICMP_HEAD					=BASE_ADDR+ETHER_ENCAP_WIDTH+VLAN_ENCAP_WIDTH+MPLS_ENCAP_WIDTH+IP_ENCAP_WIDTH;

//PARAMETERIZE THE FLOW
parameter UNIDENTIFIED_FLOW						=0;
parameter ETHER_VLAN_MPLS_IP_TCP_FLOW			=1;
parameter ETHER_VLAN_MPLS_IP_UDP_FLOW			=2;
parameter ETHER_VLAN_MPLS_IP_ICMP_FLOW			=4;
parameter ETHER_VLAN_MPLS_IP_FLOW			   =5;//
parameter ETHER_VLAN_IP_TCP_FLOW					=6;
parameter ETHER_VLAN_IP_UDP_FLOW					=7;
parameter ETHER_VLAN_IP_ICMP_FLOW				=8;
parameter ETHER_VLAN_IP_FLOW						=9;//
parameter ETHER_VLAN_ARP_FLOW						=10;
parameter ETHER_VLAN_FLOW						   =11;//
parameter ETHER_MPLS_IP_TCP_FLOW					=12;
parameter ETHER_MPLS_IP_UDP_FLOW					=13;
parameter ETHER_MPLS_IP_ICMP_FLOW				=14;
parameter ETHER_MPLS_IP_FLOW						=15;//
parameter ETHER_IP_TCP_FLOW						=16;
parameter ETHER_IP_UDP_FLOW						=17;
parameter ETHER_IP_ICMP_FLOW						=18;
parameter ETHER_IP_FLOW								=19;//
parameter ETHER_ARP_FLOW							=20;
parameter ETHER_FLOW									=21;//
parameter ERROR_FLOW									=22;

//ETHER_TYPE

parameter ETHER_TYPE_IP				=16'h0800;
parameter ETHER_TYPE_VLAN			=16'h8100;
parameter ETHER_TYPE_MPLS			=16'h8847;
parameter ETHER_TYPE_ARP			=16'h0806;

parameter VLAN_TPID_IP				=16'h0800;
parameter VLAN_TPID_VLAN			=16'h8100;
parameter VLAN_TPID_MPLS			=16'h8847;
parameter VLAN_TPID_ARP			   =16'h0806;

parameter IP_PROTOCOL_TCP			=8'h06;
parameter IP_PROTOCOL_UDP			=8'h11;
parameter IP_PROTOCOL_ICMP			=8'h01;


parameter OPENFLOW_SRC_PORT 		= 16'h6633;
parameter SWICTH_IP_ADDR    		=32'h00000000;
parameter SWICTH_MAC_ADDR			=48'h000000000000;

//parameter ADDR_WIDTH=32;

input clk;
input reset;

input glbl_program_en;

input pkt_header_ready;
output pkt_header_accept;
/*
output pkt_header_ready_accept;
input pkt_header_finish;
input pkt_header_finish_accept;


output [DPL_PKT_ADDR_WIDTH-1:0] pkt_header_addr;
input  [DPL_PKT_DATA_WIDTH-1:0] pkt_header_data;
output pkt_header_read_enable;

output reg [DPL_MATCH_FIELD_WIDTH-1:0] sdn_match_field_data;
output reg sdn_match_field_ready;
output sdn_match_field_accept;
*/
//output reg [DPL_PKT_BIT_WIDTH-1:0]pkt_header_data_buff;
output reg sdn_match_field_ready;
input [DPL_PKT_BIT_WIDTH-1:0] pkt_header_in;
output reg [DPL_PKT_BIT_WIDTH-1:0]pkt_header_data_buff;
/*
output [INGRESS_PORT_WIDTH-1:0]	sdn_ingress_port;
output [METADATA_WIDTH-1:0]		sdn_meta_data;
output [SRC_MAC_ADDR_WIDTH-1:0]	sdn_src_mac_addr;
output [DST_MAC_ADDR_WIDTH-1:0]	sdn_dst_mac_addr;
output [ETHER_TYPE_WIDTH-1:0]		sdn_ether_type;
output [VLAN_ID_WIDTH-1:0]			sdn_vlan_id;
output [VLAN_PRIORITY_WIDTH-1:0]	sdn_vlan_priority;
output [MPLS_LABEL_WIDTH-1:0]		sdn_mpls_label;
output [MPLS_FEC_WIDTH-1:0]		sdn_mpls_fec_class;
output [IP_SRC_ADDR_WIDTH-1:0]	sdn_src_ipv4_addr;
output [IP_DST_ADDR_WIDTH-1:0]	sdn_dst_ipv4_addr;
output [IP_PROTOCOL_WIDTH-1:0]	sdn_ipv4_protocol;
output [IP_TOS_WIDTH-1:0]			sdn_ipv4_tos;
output [TCP_SRC_PORT_WIDTH-1:0]	sdn_tcp_src_port;
output [TCP_DST_PORT_WIDTH-1:0]	sdn_tcp_dst_port;
*/
output reg[INGRESS_PORT_WIDTH-1:0]	OF_INGRESS_PORT;
output reg[METADATA_WIDTH-1:0]		OF_META_DATA;
output reg[SRC_MAC_ADDR_WIDTH-1:0]	OF_SRC_MAC_ADDR;
output reg[DST_MAC_ADDR_WIDTH-1:0]	OF_DST_MAC_ADDR;
output reg[ETHER_TYPE_WIDTH-1:0]		OF_ETHER_TYPE;
output reg[VLAN_ID_WIDTH-1:0]			OF_VLAN_ID;
output reg[VLAN_PRIORITY_WIDTH-1:0]	OF_VLAN_PRIORITY;
output reg[MPLS_LABEL_WIDTH-1:0]		OF_MPLS_LABEL;
output reg[MPLS_FEC_WIDTH-1:0]		OF_MPLS_FEC_CLASS;
output reg[IP_SRC_ADDR_WIDTH-1:0]	OF_SRC_IPV4_ADDR;
output reg[IP_DST_ADDR_WIDTH-1:0]	OF_DST_IPV4_ADDR;
output reg[IP_PROTOCOL_WIDTH-1:0]	OF_IP_PROTOCOL;
output reg[IP_TOS_WIDTH-1:0]			OF_IPV4_TOS;
output reg[TCP_SRC_PORT_WIDTH-1:0]	OF_TCP_SRC_PORT;
output reg[TCP_DST_PORT_WIDTH-1:0]	OF_TCP_DST_PORT;

output reg [OF_FLOW_TAG_WIDTH-1:0] of_flow_tag;
output openflow_packet_found;
output packet_to_switch_found;

output reg[ADDR_WIDTH-1:0]	OF_INGRESS_PORT_ADDR;
output reg[ADDR_WIDTH-1:0]OF_META_DATA_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_SRC_MAC_ADDR_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_DST_MAC_ADDR_ADDR;
output reg[ADDR_WIDTH-1:0] OF_ETHER_TYPE_ADDR;
output reg[ADDR_WIDTH-1:0]			OF_VLAN_ID_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_VLAN_PRIORITY_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_MPLS_LABEL_ADDR;
output reg[ADDR_WIDTH-1:0]		OF_MPLS_FEC_CLASS_ADDR;
output reg[ADDR_WIDTH-1:0]OF_SRC_IPV4_ADDR_ADDR;
output reg[ADDR_WIDTH-1:0]OF_DST_IPV4_ADDR_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_IP_PROTOCOL_ADDR;
output reg[ADDR_WIDTH-1:0]		OF_IPV4_TOS_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_TCP_SRC_PORT_ADDR;
output reg[ADDR_WIDTH-1:0]	OF_TCP_DST_PORT_ADDR;

output [DPL_MATCH_FIELD_WIDTH-1:0] OF_MATCH_FIELD_DATA;
output reg OF_FLOW_FOUND;
output reg [DPL_PKT_BIT_WIDTH-1:0] pkt_header_out;
//reg [DPL_PKT_BIT_WIDTH-1:0] pkt_header_out_buff;
/*parameter DPL_PKT_BYTE_WIDTH=64;
parameter DPL_PKT_BIT_WIDTH=512;
parameter DPL_MATCH_FIELD_WIDTH=356;
parameter DPL_PKT_ADDR_WIDTH=6;
parameter DPL_PKT_DATA_WIDTH=8;
*/
/*
assign sdn_ingress_port		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
assign sdn_meta_data			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
assign sdn_src_mac_addr    =pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
assign sdn_dst_mac_addr    =pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
assign sdn_ether_type		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];

assign sdn_vlan_id			=0;
assign sdn_vlan_priority	=0;
assign sdn_mpls_label		=0;
assign sdn_mpls_fec_class	=0;
assign sdn_src_ipv4_addr	=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
assign sdn_dst_ipv4_addr	=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
assign sdn_ipv4_protocol	=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
assign sdn_ipv4_tos			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
assign sdn_tcp_src_port		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
assign sdn_tcp_dst_port  	=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
*/
reg pkt_header_accept;
reg pkt_header_data_valid;


wire [ETHER_TYPE_WIDTH-1:0] ether_type;
wire [VLAN_TPID_WIDTH-1:0]	 ether_vlan_flow_ether_type;
wire [IP_PROTOCOL_WIDTH-1:0] ether_ip_flow_ip_protocol;
wire [IP_PROTOCOL_WIDTH-1:0] ether_vlan_ip_flow_ip_protocol;
wire [IP_PROTOCOL_WIDTH-1:0] ether_mpls_ip_flow_ip_protocol;
wire [IP_PROTOCOL_WIDTH-1:0] ether_vlan_mpls_ip_flow_ip_protocol;

assign ether_type										=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
assign ether_vlan_flow_ether_type				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_FLOW_VLAN_HEAD+32)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_FLOW_VLAN_HEAD+32+ETHER_TYPE_WIDTH))];
assign ether_ip_flow_ip_protocol					=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
assign ether_vlan_ip_flow_ip_protocol			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
assign ether_mpls_ip_flow_ip_protocol			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
assign ether_vlan_mpls_ip_flow_ip_protocol	=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];

assign OF_MATCH_FIELD_DATA={  OF_INGRESS_PORT,OF_META_DATA,OF_DST_MAC_ADDR, OF_SRC_MAC_ADDR, OF_ETHER_TYPE, OF_VLAN_ID, OF_VLAN_PRIORITY, OF_MPLS_LABEL, OF_MPLS_FEC_CLASS, OF_SRC_IPV4_ADDR, OF_DST_IPV4_ADDR, OF_IP_PROTOCOL, OF_IPV4_TOS, OF_TCP_SRC_PORT, OF_TCP_DST_PORT};
//Parameter of The Header Fileds
initial begin
pkt_header_data_valid<=1'b0;
end


always@(posedge clk)begin
 //$display("%g %b",$time,clk);
   if(!reset)begin
	if(!glbl_program_en)begin
       if(pkt_header_ready)begin
             pkt_header_data_buff<=pkt_header_in;
               pkt_header_accept<=1'b1;
			      pkt_header_data_valid<=1'b1;
			
      end
      else begin
         pkt_header_data_buff<=pkt_header_data_buff;
         pkt_header_data_valid<=0;
          pkt_header_accept<=1'b0;
      end	//
	  end//GLBL PROG
   end 
	else begin
			pkt_header_data_buff<=0;
         pkt_header_accept<=1'b0;
			pkt_header_data_valid<=1'b0;
	end
end

always@(posedge clk)begin
if(!reset)begin
  if(!glbl_program_en)begin
  //$display("%g ether_type: %x \n ether_vlan_flow_ether_type: %x \n ether_ip_flow_ip_protocol: %x \n ether_vlan_ip_flow_ip_protocol: %x \n  ether_mpls_ip_flow_ip_protocol: %x\n ether_vlan_mpls_ip_flow_ip_protocol: %x\n",$time,ether_type,ether_vlan_flow_ether_type,ether_ip_flow_ip_protocol,ether_vlan_ip_flow_ip_protocol,ether_mpls_ip_flow_ip_protocol,ether_vlan_mpls_ip_flow_ip_protocol);
  	if(pkt_header_data_valid)begin
			pkt_header_out<=pkt_header_data_buff;
				if(ether_type==ETHER_TYPE_VLAN )begin 
			      if(ether_vlan_flow_ether_type==ETHER_TYPE_MPLS)begin
							if(ether_vlan_mpls_ip_flow_ip_protocol==IP_PROTOCOL_TCP)begin
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
						      
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1;

								sdn_match_field_ready=1'b1;
								OF_FLOW_FOUND=1'b1;
								of_flow_tag<=ETHER_VLAN_MPLS_IP_TCP_FLOW;
								
								/*if(OF_TCP_SRC_PORT ==OPENFLOW_SRC_PORT )begin
								      openflow_packet_found=1;
								end
								else begin
								     openflow_packet_found=0;
								end
								
								if(OF_DST_IPV4_ADDR == SWICTH_IP_ADDR)begin
								     packet_to_switch_found=1;
								end
								else begin
								    packet_to_switch_found=0;
								end*/
								//$display("FLOW: ETHER_VLAN_MPLS_TCP\n");
						end
							if(ether_vlan_mpls_ip_flow_ip_protocol==IP_PROTOCOL_UDP)begin
									
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1;
									 
									 
									 sdn_match_field_ready=1'b1;
								     OF_FLOW_FOUND=1'b1;
									  of_flow_tag<=ETHER_VLAN_MPLS_IP_UDP_FLOW;
									 //$display("FLOW: ETHER_VLAN_MPLS_UDP\n");
									/*if(OF_UDP_SRC_PORT ==OPENFLOW_SRC_PORT )begin
								      openflow_packet_found=1;
									end
									else begin
								     openflow_packet_found=0;
									end
								
									if(OF_DST_IPV4_ADDR == SWICTH_IP_ADDR)begin
								     packet_to_switch_found=1;
									end
									else begin
								    packet_to_switch_found=0;
									end*/
									 
									 
							end
							if(ether_vlan_mpls_ip_flow_ip_protocol==IP_PROTOCOL_ICMP)begin
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;									
									
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_VLAN_MPLS_IP_ICMP_FLOW;
									// $display("FLOW: ETHER_VLAN_MPLS_ICMP\n");
									/*
									openflow_packet_found=0;									
								
									if(OF_DST_IPV4_ADDR == SWICTH_IP_ADDR)begin
								     packet_to_switch_found=1;
									end
									else begin
								    packet_to_switch_found=0;
									end*/
							end
							else begin
									
									OF_INGRESS_PORT	=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_VLAN_MPLS_IP_FLOW;
									
								   /*openflow_packet_found=0;
									
									if(OF_DST_IPV4_ADDR == SWICTH_IP_ADDR)begin
								     packet_to_switch_found=1;
									end
									else begin
								    packet_to_switch_found=0;
									end*/
									
							     //$display("ERROR: UNIDENTIFIED FLOW - ETHER_VLAN_MPLS_IP?\n");
							end					     
					end
					else if(ether_vlan_flow_ether_type==ETHER_TYPE_IP)begin
							if(ether_vlan_ip_flow_ip_protocol==IP_PROTOCOL_TCP)begin
							      OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
							       
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1;
									
									 
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_VLAN_IP_TCP_FLOW;
									/*
									if(OF_TCP_SRC_PORT ==OPENFLOW_SRC_PORT )begin
								      openflow_packet_found=1;
									end
									else begin
								     openflow_packet_found=0;
									end
								
									if(OF_DST_IPV4_ADDR == SWICTH_IP_ADDR)begin
								     packet_to_switch_found=1;
									end
									else begin
								    packet_to_switch_found=0;
									end*/
									// $display("FLOW: ETHER_VLAN_IP_TCP\n");
							end
							if(ether_vlan_ip_flow_ip_protocol==IP_PROTOCOL_UDP)begin
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
									 
									 
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1;
									 
									 
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_VLAN_IP_UDP_FLOW;
									 $display("FLOW: ETHER_VLAN_IP_UDP\n");
							end
							if(ether_vlan_ip_flow_ip_protocol==IP_PROTOCOL_ICMP)begin
							    
								   OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									
									 
									 sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_VLAN_IP_ICMP_FLOW;
									 $display("FLOW: ETHER_VLAN_IP_ICMP\n");
						
							end
							else begin
							    $display("ERROR: UNIDENTIFIED FLOW - ETHER_VLAN_IP?\n");
								   /*OF_INGRESS_PORT		=0;
									OF_META_DATA			=0;
									OF_DST_MAC_ADDR		=0;
									OF_SRC_MAC_ADDR		=0;
									OF_ETHER_TYPE			=0;
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=0;
									OF_DST_IPV4_ADDR		=0;
									OF_IP_PROTOCOL			=0;
									OF_IPV4_TOS				=0;
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									
									OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0; */
									
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;									
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_VLAN_IP_FLOW;
							end							
					end
					
					else if(ether_vlan_flow_ether_type==ETHER_TYPE_ARP)begin
					     //YET TO IMPLEMENT
						      	OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=0;
									OF_DST_IPV4_ADDR		=0;
									OF_IP_PROTOCOL			=0;
									OF_IPV4_TOS				=0;
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;	
									
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_VLAN_ARP_FLOW;
									 $display("FLOW: ETHER_VLAN_ARP\n");
					end
					else begin
					$display("ERROR: UNIDENTIFIED FLOW - ETHER_VLAN?\n");
					            /*OF_INGRESS_PORT		=0;
									OF_META_DATA			=0;
									OF_DST_MAC_ADDR		=0;
									OF_SRC_MAC_ADDR		=0;
									OF_ETHER_TYPE			=0;
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=0;
									OF_DST_IPV4_ADDR		=0;
									OF_IP_PROTOCOL			=0;
									OF_IPV4_TOS				=0;
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;									
									
									
									OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
									*/
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET+VLAN_ID_WIDTH))];
									OF_VLAN_PRIORITY		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET+VLAN_PRIORITY_WIDTH))];
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=0;
									OF_DST_IPV4_ADDR		=0;
									OF_IP_PROTOCOL			=0;
									OF_IPV4_TOS				=0;
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;	
									
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_ID_OFFSET)-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_VLAN_ARP_FLOW_VLAN_HEAD+VLAN_PRIORITY_OFFSET)-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;

									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;	
										of_flow_tag<=ETHER_VLAN_FLOW;
									
					end
					
			end//END ETHER_TYPE_MPLS
			else if(ether_type==ETHER_TYPE_MPLS)begin
					if(ether_mpls_ip_flow_ip_protocol==IP_PROTOCOL_TCP)begin
							      OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
								
								
								   OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1;
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_MPLS_IP_TCP_FLOW;
								$display("FLOW: ETHER_MPLS_IP_TCP\n");
					
					end
					else if(ether_mpls_ip_flow_ip_protocol==IP_PROTOCOL_UDP)begin
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
									OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
					      	
								   OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1;
								
								
								
								sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_MPLS_IP_UDP_FLOW;
							$display("FLOW: ETHER_MPLS_IP_UDP\n");
					end
					else if(ether_mpls_ip_flow_ip_protocol==IP_PROTOCOL_ICMP)begin
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									
									 OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									
									
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_MPLS_IP_ICMP_FLOW;
									$display("FLOW: ETHER_MPLS_IP_ICMP\n");
					
					end
					else begin
					            $display("ERROR: UNIDENTIFIED FLOW - ETHER_MPLS?\n");
									/*OF_INGRESS_PORT		=0;
									OF_META_DATA			=0;
									OF_DST_MAC_ADDR		=0;
									OF_SRC_MAC_ADDR		=0;
									OF_ETHER_TYPE			=0;
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=0;
									OF_MPLS_FEC_CLASS		=0;
									OF_SRC_IPV4_ADDR		=0;
									OF_DST_IPV4_ADDR		=0;
									OF_IP_PROTOCOL			=0;
									OF_IPV4_TOS				=0;
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
									*/
									
									OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
									OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
									OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
									OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
									OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
									OF_VLAN_ID				=0;
									OF_VLAN_PRIORITY		=0;
									OF_MPLS_LABEL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET+MPLS_LABEL_WIDTH))];
									OF_MPLS_FEC_CLASS		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET+MPLS_FEC_CLASS_WIDTH))];
									OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
									OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
									OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
									OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
									OF_TCP_SRC_PORT		=0;
									OF_TCP_DST_PORT		=0;
									
									
									OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_LABEL_OFFSET)-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_MPLS_HEAD+MPLS_FEC_CLASS_OFFSET)-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_MPLS_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									
									sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_MPLS_IP_FLOW;
					
					end
			end//END ETHER_TYPE_MPLS
			
			else if(ether_type==ETHER_TYPE_IP)begin
					if(ether_ip_flow_ip_protocol==IP_PROTOCOL_TCP)begin
					      
						OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
						OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
						OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
						OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
						OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET+TCP_SRC_PORT_WIDTH))];
						OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET+TCP_DST_PORT_WIDTH))];
						
						
							      OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_TCP_FLOW_TCP_HEAD+TCP_DST_PORT_OFFSET)-1;
									
							     sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
									of_flow_tag<=ETHER_IP_TCP_FLOW;
						$display("FLOW: ETHER_IP_TCP\n");
					end
					else if(ether_ip_flow_ip_protocol==IP_PROTOCOL_UDP)begin
					     
						OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
						OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
						OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
						OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
						OF_TCP_SRC_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET+UDP_SRC_PORT_WIDTH))];
						OF_TCP_DST_PORT		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET+UDP_DST_PORT_WIDTH))];
						
							      OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_SRC_PORT_OFFSET)-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_UDP_FLOW_UDP_HEAD+UDP_DST_PORT_OFFSET)-1;
						
							sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_IP_UDP_FLOW;
						$display("FLOW: ETHER_IP_UDP\n");
					end
					else if(ether_ip_flow_ip_protocol==IP_PROTOCOL_ICMP)begin
					   OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
						OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
						OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
						OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
							      OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
							
							sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_IP_ICMP_FLOW;
						$display("FLOW: ETHER_IP_ICMP\n");
					end
					else begin
					    $display("ERROR: UNIDENTIFIED FLOW - ETHER_IP?\n");
				      /* OF_INGRESS_PORT		=0;
						OF_META_DATA			=0;
						OF_DST_MAC_ADDR		=0;
						OF_SRC_MAC_ADDR		=0;
						OF_ETHER_TYPE			=0;
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
					         	OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
									*/
									  OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET+IP_SRC_ADDR_WIDTH))];
						OF_DST_IPV4_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET+IP_DST_ADDR_WIDTH))];
						OF_IP_PROTOCOL			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET+IP_PROTOCOL_WIDTH))];
						OF_IPV4_TOS				=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(ETHER_IP_FLOW_IP_HEAD+IP_TOS_OFFSET+IP_TOS_WIDTH))];
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
							      OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_SRC_ADDR_OFFSET)-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_DST_ADDR_OFFSET)-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_PROTOCOL_OFFSET)-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-(ETHER_IP_ICMP_FLOW_IP_HEAD+IP_TOS_OFFSET)-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
						
							sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_IP_FLOW;
					end			
			end//END ETHER_TYPE_IP
			else if (ether_type==ETHER_TYPE_ARP)begin
					   OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
						         OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
						
							sdn_match_field_ready=1'b1;
								   OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_ARP_FLOW;
						$display("FLOW: ETHER_ARP\n");
					
			end
			else begin
			    $display("ERROR: UNIDENTIFIED FLOW - ETHER? \n");
				      /*OF_INGRESS_PORT		=0;
						OF_META_DATA			=0;
						OF_DST_MAC_ADDR		=0;
						OF_SRC_MAC_ADDR		=0;
						OF_ETHER_TYPE			=0;
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
						         OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
									
									*/
									
									 OF_INGRESS_PORT		=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-ROOT_ADDR-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+INGRESS_PORT_OFFSET+INGRESS_PORT_WIDTH))];
						OF_META_DATA			=pkt_header_data_buff[DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1:(DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET+METADATA_WIDTH))];
						OF_DST_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET+DST_MAC_ADDR_WIDTH))];
						OF_SRC_MAC_ADDR		=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET+SRC_MAC_ADDR_WIDTH))];
						OF_ETHER_TYPE			=pkt_header_data_buff[(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1):(DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET+ETHER_TYPE_WIDTH))];
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
						         OF_INGRESS_PORT_ADDR		=DPL_PKT_BIT_WIDTH-ROOT_ADDR-1;
									OF_META_DATA_ADDR			=DPL_PKT_BIT_WIDTH-(ROOT_ADDR+METADATA_OFFSET)-1;
									OF_DST_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_DST_OFFSET)-1;
									OF_SRC_MAC_ADDR_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+MAC_SRC_OFFSET)-1;
									OF_ETHER_TYPE_ADDR		=DPL_PKT_BIT_WIDTH-(BASE_ADDR+ETHER_TYPE_OFFSET)-1;
									OF_VLAN_ID_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_VLAN_PRIORITY_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_LABEL_ADDR      =DPL_PKT_BIT_WIDTH-1;
									OF_MPLS_FEC_CLASS_ADDR  =DPL_PKT_BIT_WIDTH-1;
									OF_SRC_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_DST_IPV4_ADDR_ADDR	=DPL_PKT_BIT_WIDTH-1;
									OF_IP_PROTOCOL_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_IPV4_TOS_ADDR			=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_SRC_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
									OF_TCP_DST_PORT_ADDR		=DPL_PKT_BIT_WIDTH-1;
						
							       sdn_match_field_ready=1'b1;
								    OF_FLOW_FOUND=1'b1;
										of_flow_tag<=ETHER_FLOW;			    
			end				
	   end//VALID	
		else begin
						OF_INGRESS_PORT		=0;
						OF_META_DATA			=0;
						OF_DST_MAC_ADDR		=0;
						OF_SRC_MAC_ADDR		=0;
						OF_ETHER_TYPE			=0;
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
					         	OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
		               
		                       sdn_match_field_ready=1'b0;
								   OF_FLOW_FOUND=1'b0;
		end
	 end//GLBL PROGRAM	
   end//RESET	
	else begin
				OF_INGRESS_PORT		=0;
						OF_META_DATA			=0;
						OF_DST_MAC_ADDR		=0;
						OF_SRC_MAC_ADDR		=0;
						OF_ETHER_TYPE			=0;
						OF_VLAN_ID				=0;
						OF_VLAN_PRIORITY		=0;
						OF_MPLS_LABEL			=0;
						OF_MPLS_FEC_CLASS		=0;
						OF_SRC_IPV4_ADDR		=0;
						OF_DST_IPV4_ADDR		=0;
						OF_IP_PROTOCOL			=0;
						OF_IPV4_TOS				=0;
						OF_TCP_SRC_PORT		=0;
						OF_TCP_DST_PORT		=0;
						
					         	OF_INGRESS_PORT_ADDR		=0;
									OF_META_DATA_ADDR			=0;
									OF_DST_MAC_ADDR_ADDR		=0;
									OF_SRC_MAC_ADDR_ADDR		=0;
									OF_ETHER_TYPE_ADDR		=0;
									OF_VLAN_ID_ADDR			=0;
									OF_VLAN_PRIORITY_ADDR	=0;
									OF_MPLS_LABEL_ADDR      =0;
									OF_MPLS_FEC_CLASS_ADDR  =0;
									OF_SRC_IPV4_ADDR_ADDR	=0;
									OF_DST_IPV4_ADDR_ADDR	=0;
									OF_IP_PROTOCOL_ADDR		=0;
									OF_IPV4_TOS_ADDR			=0;
									OF_TCP_SRC_PORT_ADDR		=0;
									OF_TCP_DST_PORT_ADDR		=0;
		               
		                       sdn_match_field_ready=1'b0;
								   OF_FLOW_FOUND=1'b0;
	
	end
	
	
end

/*
always@(posedge clk) begin
if(!reset)begin
  if(pkt_header_data_valid)begin
    sdn_match_field_data<=pkt_header_data_buff[355:0];
	 pkt_header_data_valid<=1'b0;
	end
end

end
endmodule

*/

endmodule
