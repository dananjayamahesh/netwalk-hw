`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:24:53 01/11/2016 
// Design Name: 
// Module Name:    netwalk_encoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module netwalk_encoder
#(parameter ENCODER_OUT_WIDTH=6)
(
clk,
reset,
encoder_in,
encoder_out
);
parameter ENCODER_IN_WIDTH=1<<ENCODER_OUT_WIDTH;
input clk;
input reset;
input [ENCODER_IN_WIDTH-1:0]encoder_in;
output reg[ENCODER_OUT_WIDTH-1:0]encoder_out;

reg[ENCODER_OUT_WIDTH-1:0] map[0:ENCODER_IN_WIDTH-1];
reg map_set;
integer i;
integer j;

always@(*)begin
  if(!reset)begin
       case(encoder_in)
			64'b0000000000000000000000000000000000000000000000000000000000000001: encoder_out<=6'b000000;
			64'b0000000000000000000000000000000000000000000000000000000000000010: encoder_out<=6'b000001;
			64'b0000000000000000000000000000000000000000000000000000000000000100: encoder_out<=6'b000010;
			64'b0000000000000000000000000000000000000000000000000000000000001000: encoder_out<=6'b000011;
			64'b0000000000000000000000000000000000000000000000000000000000010000: encoder_out<=6'b000100;
			64'b0000000000000000000000000000000000000000000000000000000000100000: encoder_out<=6'b000101;
			64'b0000000000000000000000000000000000000000000000000000000001000000: encoder_out<=6'b000110;
			64'b0000000000000000000000000000000000000000000000000000000010000000: encoder_out<=6'b000111;
			64'b0000000000000000000000000000000000000000000000000000000100000000: encoder_out<=6'b001000;
			64'b0000000000000000000000000000000000000000000000000000001000000000: encoder_out<=6'b001001;
			64'b0000000000000000000000000000000000000000000000000000010000000000: encoder_out<=6'b001010;
			64'b0000000000000000000000000000000000000000000000000000100000000000: encoder_out<=6'b001011;
			64'b0000000000000000000000000000000000000000000000000001000000000000: encoder_out<=6'b001100;
			64'b0000000000000000000000000000000000000000000000000010000000000000: encoder_out<=6'b001101;
			64'b0000000000000000000000000000000000000000000000000100000000000000: encoder_out<=6'b001110;
			64'b0000000000000000000000000000000000000000000000001000000000000000: encoder_out<=6'b001111;
			64'b0000000000000000000000000000000000000000000000010000000000000000: encoder_out<=6'b010000;
			64'b0000000000000000000000000000000000000000000000100000000000000000: encoder_out<=6'b010001;
			64'b0000000000000000000000000000000000000000000001000000000000000000: encoder_out<=6'b010010;
			64'b0000000000000000000000000000000000000000000010000000000000000000: encoder_out<=6'b010011;
			64'b0000000000000000000000000000000000000000000100000000000000000000: encoder_out<=6'b010100;
			64'b0000000000000000000000000000000000000000001000000000000000000000: encoder_out<=6'b010101;
			64'b0000000000000000000000000000000000000000010000000000000000000000: encoder_out<=6'b010110;
			64'b0000000000000000000000000000000000000000100000000000000000000000: encoder_out<=6'b010111;
			64'b0000000000000000000000000000000000000001000000000000000000000000: encoder_out<=6'b011000;
			64'b0000000000000000000000000000000000000010000000000000000000000000: encoder_out<=6'b011001;
			64'b0000000000000000000000000000000000000100000000000000000000000000: encoder_out<=6'b011010;
			64'b0000000000000000000000000000000000001000000000000000000000000000: encoder_out<=6'b011011;
			64'b0000000000000000000000000000000000010000000000000000000000000000: encoder_out<=6'b011100;
			64'b0000000000000000000000000000000000100000000000000000000000000000: encoder_out<=6'b011101;
			64'b0000000000000000000000000000000001000000000000000000000000000000: encoder_out<=6'b011110;
			64'b0000000000000000000000000000000010000000000000000000000000000000: encoder_out<=6'b011111;
			64'b0000000000000000000000000000000100000000000000000000000000000000: encoder_out<=6'b100000;
			64'b0000000000000000000000000000001000000000000000000000000000000000: encoder_out<=6'b100001;
			64'b0000000000000000000000000000010000000000000000000000000000000000: encoder_out<=6'b100010;
			64'b0000000000000000000000000000100000000000000000000000000000000000: encoder_out<=6'b100011;
			64'b0000000000000000000000000001000000000000000000000000000000000000: encoder_out<=6'b100100;
			64'b0000000000000000000000000010000000000000000000000000000000000000: encoder_out<=6'b100101;
			64'b0000000000000000000000000100000000000000000000000000000000000000: encoder_out<=6'b100110;
			64'b0000000000000000000000001000000000000000000000000000000000000000: encoder_out<=6'b100111;
			64'b0000000000000000000000010000000000000000000000000000000000000000: encoder_out<=6'b101000;
			64'b0000000000000000000000100000000000000000000000000000000000000000: encoder_out<=6'b101001;
			64'b0000000000000000000001000000000000000000000000000000000000000000: encoder_out<=6'b101010;
			64'b0000000000000000000010000000000000000000000000000000000000000000: encoder_out<=6'b101011;
			64'b0000000000000000000100000000000000000000000000000000000000000000: encoder_out<=6'b101100;
			64'b0000000000000000001000000000000000000000000000000000000000000000: encoder_out<=6'b101101;
			64'b0000000000000000010000000000000000000000000000000000000000000000: encoder_out<=6'b101110;
			64'b0000000000000000100000000000000000000000000000000000000000000000: encoder_out<=6'b101111;
			64'b0000000000000001000000000000000000000000000000000000000000000000: encoder_out<=6'b110000;
			64'b0000000000000010000000000000000000000000000000000000000000000000: encoder_out<=6'b110001;
			64'b0000000000000100000000000000000000000000000000000000000000000000: encoder_out<=6'b110010;
			64'b0000000000001000000000000000000000000000000000000000000000000000: encoder_out<=6'b110011;
			64'b0000000000010000000000000000000000000000000000000000000000000000: encoder_out<=6'b110100;
			64'b0000000000100000000000000000000000000000000000000000000000000000: encoder_out<=6'b110101;
			64'b0000000001000000000000000000000000000000000000000000000000000000: encoder_out<=6'b110110;
			64'b0000000010000000000000000000000000000000000000000000000000000000: encoder_out<=6'b110111;
			64'b0000000100000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111000;
			64'b0000001000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111001;
			64'b0000010000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111010;
			64'b0000100000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111011;
			64'b0001000000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111100;
			64'b0010000000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111101;
			64'b0100000000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111110;
			64'b1000000000000000000000000000000000000000000000000000000000000000: encoder_out<=6'b111111;
			default: encoder_out<=6'b111111;

	 endcase
  end
    
  else begin
  encoder_out<=6'b000000;
  end
end


/*
always@(posedge clk) begin
   if(encoder_enable)begin
	  if(!reset)begin
			if(!map_set)begin
		      for(j=0;j<ENCODER_IN_WIDTH;j=j+1)begin
				     map[j] <= j;
				end	
           map_set<=1;				
			end	
			else begin
		      map_set<=1;
			end 
	  end
	  else begin
	     map_set<=0;
	  end  
	end  
	else begin
	     map_set<=0;	  
	 end  
end
	  
always@(encoder_in)begin
  if(encoder_enable)begin
		if(!reset)begin
		   for(i=0;i<ENCODER_IN_WIDTH;i=i+1)begin
			       if(encoder_in[i]==1'b1)begin
					        encoder_out <= map[i];					 
					 end
		 	end
		end
		else begin
          encoder_out<=0;
		end		
	end
   else begin
     encoder_out<=0;
	end	
end
*/

endmodule

